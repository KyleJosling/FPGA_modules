// localparam reg [COEFF_WIDTH-1:0] coeff_array[0:127] = '{128{18'h00020}};                                        
localparam reg [COEFF_WIDTH-1:0] coeff_array[0:127] = '{18'h3FBFB,
                                                      18'h3F61D,
                                                      18'h3F5F4,
                                                      18'h3FBC5,
                                                      18'h0044D,
                                                      18'h00A90,
                                                      18'h00ABF,
                                                      18'h00487,
                                                      18'h3FB64,
                                                      18'h3F4AA,
                                                      18'h3F473,
                                                      18'h3FB20,
                                                      18'h004F8,
                                                      18'h00C3C,
                                                      18'h00C7C,
                                                      18'h00547,
                                                      18'h3FA9D,
                                                      18'h3F2B6,
                                                      18'h3F26B,
                                                      18'h3FA40,
                                                      18'h005E2,
                                                      18'h00E8A,
                                                      18'h00EE4,
                                                      18'h00652,
                                                      18'h3F985,
                                                      18'h3EFF3,
                                                      18'h3EF85,
                                                      18'h3F8FD,
                                                      18'h00736,
                                                      18'h011E9,
                                                      18'h01272,
                                                      18'h007E0,
                                                      18'h3F7E0,
                                                      18'h3EBBD,
                                                      18'h3EB0D,
                                                      18'h3F705,
                                                      18'h0094F,
                                                      18'h01752,
                                                      18'h0183C,
                                                      18'h00A72,
                                                      18'h3F51C,
                                                      18'h3E489,
                                                      18'h3E342,
                                                      18'h3F384,
                                                      18'h00D20,
                                                      18'h02168,
                                                      18'h02350,
                                                      18'h00F83,
                                                      18'h3EF7C,
                                                      18'h3D561,
                                                      18'h3D239,
                                                      18'h3EB86,
                                                      18'h01642,
                                                      18'h03ADC,
                                                      18'h0410E,
                                                      18'h01E1E,
                                                      18'h3DDDE,
                                                      18'h3A0EB,
                                                      18'h38FA2,
                                                      18'h3C71D,
                                                      18'h04924,
                                                      18'h0F736,
                                                      18'h19C05,
                                                      18'h1FFFF,
                                                      18'h1FFFF,
                                                      18'h19C05,
                                                      18'h0F736,
                                                      18'h04924,
                                                      18'h3C71D,
                                                      18'h38FA2,
                                                      18'h3A0EB,
                                                      18'h3DDDE,
                                                      18'h01E1E,
                                                      18'h0410E,
                                                      18'h03ADC,
                                                      18'h01642,
                                                      18'h3EB86,
                                                      18'h3D239,
                                                      18'h3D561,
                                                      18'h3EF7C,
                                                      18'h00F83,
                                                      18'h02350,
                                                      18'h02168,
                                                      18'h00D20,
                                                      18'h3F384,
                                                      18'h3E342,
                                                      18'h3E489,
                                                      18'h3F51C,
                                                      18'h00A72,
                                                      18'h0183C,
                                                      18'h01752,
                                                      18'h0094F,
                                                      18'h3F705,
                                                      18'h3EB0D,
                                                      18'h3EBBD,
                                                      18'h3F7E0,
                                                      18'h007E0,
                                                      18'h01272,
                                                      18'h011E9,
                                                      18'h00736,
                                                      18'h3F8FD,
                                                      18'h3EF85,
                                                      18'h3EFF3,
                                                      18'h3F985,
                                                      18'h00652,
                                                      18'h00EE4,
                                                      18'h00E8A,
                                                      18'h005E2,
                                                      18'h3FA40,
                                                      18'h3F26B,
                                                      18'h3F2B6,
                                                      18'h3FA9D,
                                                      18'h00547,
                                                      18'h00C7C,
                                                      18'h00C3C,
                                                      18'h004F8,
                                                      18'h3FB20,
                                                      18'h3F473,
                                                      18'h3F4AA,
                                                      18'h3FB64,
                                                      18'h00487,
                                                      18'h00ABF,
                                                      18'h00A90,
                                                      18'h0044D,
                                                      18'h3FBC5,
                                                      18'h3F5F4,
                                                      18'h3F61D,
                                                      18'h3FBF8};
